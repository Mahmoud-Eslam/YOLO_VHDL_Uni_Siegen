library IEEE;
use IEEE.std_logic_1164.ALL;
use IEEE.std_logic_arith.ALL;
use IEEE.math_real.ALL;

package conv_package is 
    type integer_1d_vector is array(integer range <>) of integer;
    type float_1d_vector is array(Natural range <>) of real;
    
    type integer_2d_vector is array(integer range <>, integer range <>) of integer;
    type float_2d_vector is array(Natural range <>, Natural range <>) of real;
    
    type integer_3d_vector is array(integer range <>, integer range <>, integer range <>) of integer;
    type float_3d_vector is array(Natural range <>, Natural range <>, Natural range <>) of real;
    
    type integer_4d_vector is array(integer range <>, integer range <>, integer range <>, integer range <>) of integer;
    type float_4d_vector is array(Natural range <>, Natural range <>, Natural range <>, Natural range <>) of real;
end;    	

library IEEE;
use IEEE.std_logic_1164.ALL;
use IEEE.std_logic_arith.ALL;
use IEEE.math_real.ALL;

library work;
use work.conv_package.all;

entity YOLO_VHDL_Source is 
    generic(            
            pooled_height :integer := 15;
            pooled_width  :integer := 15;
            i_filters     :integer := 16;
            stride        :integer := 2
            );
    port(
        CLK : in std_logic;
        reset : in std_logic;
        new_img : out float_3d_vector (0 to (pooled_height - 1), 0 to (pooled_width - 1), 0 to (i_filters - 1)) := (others => (others => (others => 0.0)))
        );       
end YOLO_VHDL_Source;

architecture Behavioral of YOLO_VHDL_Source is  
 
constant i_height  :integer := 32; 
constant i_width   :integer := 32;
constant i_depth   :integer := 3; 
 
constant img : float_3d_vector :=
    (
    ((0.8619490974451727, 6.669539947472779, 7.962096925143088), (4.928269279891456, 7.509230450500263, 7.5805488465059465), (8.76414636327273, 2.509301100106194, 1.3493890300535571), (8.200251891197368, 5.966745801655534, 7.680102152799526), (2.0552140419517126, 8.671417205339004, 3.169678449947585), (2.963212432601121, 6.532063992562963, 8.412180238497827), (7.790390118369049, 5.022881515193983, 1.346444711063245), (3.9410427877245793, 5.645238770366055, 3.8371263271413234), (4.156071526671676, 2.9498920054823063, 9.934693510317645), (2.894852004692302, 1.3770149990694214, 5.277773894756842), (2.0902486554260067, 1.4118559244493056, 9.408311888411426), (3.6019829035614492, 3.9368926772480464, 7.119552891797678), (5.179680159737602, 7.306112305603265, 0.5491565240270646), (5.588299765659453, 1.7677475882892313, 9.581706752168571), (6.754027543418032, 9.487468383177278, 9.015613183608451), (0.6741380958239873, 7.771434476471554, 9.497761615198172), (2.450284288129688, 8.554991826711277, 1.379162842516396), (2.067195918596947, 5.193354608772101, 7.009781844436099), (2.0499044241676865, 6.747512949002521, 0.34290735858084287), (0.8206640638035867, 8.9180882669109, 1.1413528319957411), (2.6652282911639236, 6.177629764067244, 9.900312797302256), (8.632785426045954, 0.028979754922677792, 0.5918027450514185), (5.483393986562427, 7.157783777954135, 2.9818115623016483), (0.5439779066201111, 4.487425510442582, 0.6188275128572529), (1.2405502316922368, 2.52221594903292, 5.184389103277251), (1.6782975883643292, 1.6552578136198193, 2.8202279035451716), (1.676966863496887, 3.0458634661248585, 6.964632649852234), (1.275339036104145, 1.2907723274548333, 8.844547588064911), (2.7202201087152265, 3.0201126964593783, 7.894539362120028), (6.695096577964889, 2.453300380192631, 9.22044177933206), (1.7314440965186295, 3.6543973894094317, 5.183905926250313), (6.5581830805192105, 5.711929275132329, 0.21580211673071892)),
    ((9.86898446245713, 6.031441191291273, 9.694121669957587), (7.551685330938128, 4.052196305427303, 7.80458820849508), (7.1317072004986946, 7.149311800418584, 2.080473105864055), (7.37180791031135, 7.8869822719193206, 5.156421892620598), (4.545498066344496, 7.462095614890042, 1.9076243836820006), (4.348284298289727, 6.259051059058081, 1.6305730520575734), (3.3417623389797892, 3.7129122189118102, 2.883094804342762), (3.171693046979638, 6.503078768329677, 1.7817202719823955), (5.768192819927695, 2.9184149446777408, 0.5324131986380642), (0.9590580639654245, 4.001675075989723, 3.1278357031364665), (6.771957297831726, 1.320327492958503, 4.8690630163245725), (4.265064158576999, 6.685214068490044, 2.310043705400413), (6.1804633839255905, 2.326507485706979, 4.591473572157065), (1.416899741979668, 9.731925059915298, 5.7980093789119325), (0.8698048593993102, 0.21331464836096048, 5.830782454096479), (8.974937217950545, 3.350790076197204, 7.382192449536989), (3.274278235819433, 1.1082402318690132, 1.1474321616520333), (3.892156350695126, 5.9156099696225715, 1.2056344548884568), (9.047784701725883, 0.8484586378625036, 9.50141853731158), (2.877562302642515, 7.8745171518207115, 1.2733511331989167), (5.920396084928758, 6.615921789676573, 0.39288145833782706), (3.741023605246747, 2.5314966417172324, 6.4155581719844275), (5.278566529091481, 2.1820962680493547, 9.730596389232115), (0.7122517540480056, 0.8843186998595476, 5.659908674350154), (8.465923180410815, 0.6983917349223523, 7.964905053497301), (2.068144035919639, 2.7197422352456146, 7.387020511646584), (4.261224710833198, 6.844859155375815, 6.731275421957054), (4.403310777615712, 8.706668093562264, 4.806545968810692), (7.959013234625171, 2.1547062102728507, 7.182252091011504), (6.823758828540569, 0.7264771460510255, 9.249724434815336), (7.906079037249777, 2.7968531535599817, 9.41331986809834), (6.5791730436307425, 1.123985361545109, 0.6897624299509608)),
    ((3.347615336436264, 7.848871556679172, 4.083756574703708), (7.053561438031655, 0.42559227483635054, 3.692114103565971), (5.5901404604589375, 5.682446729469968, 4.191510708980779), (1.3912419299803158, 6.199362194365614, 0.38579777285881467), (3.206103334580115, 9.480149525022114, 3.5722922138606594), (8.824858741139685, 2.8002091335853354, 3.9987101521013457), (8.96363989444304, 1.270088764736056, 5.340964140779025), (2.8933026019399866, 0.8371989017813342, 3.8529426308413814), (4.774088108177694, 2.049529240852992, 5.762721992897807), (1.2026808790118704, 3.4597820803794677, 8.60215703683648), (7.102892664049114, 4.676490572738468, 0.39178897632646037), (6.500424411841976, 4.075995762042308, 8.795863362700887), (4.5032434445337755, 9.2939634808245, 0.4645229704362652), (6.523759186773671, 7.025740591526351, 9.277380116676051), (7.578929699451406, 0.7986030787386067, 1.5033093086013916), (0.4691108330751004, 3.400231242421813, 2.171329971139576), (0.13912597970602847, 9.470109756290256, 9.960951330361805), (0.3546341804414932, 5.7442973680239975, 1.6094267751653635), (6.806357249218821, 0.6860107164250051, 6.340337098305422), (2.9010739774957317, 7.888334700056792, 4.795816170653016), (1.565005766849118, 0.5817352194212444, 6.123869353893941), (3.0092409338034987, 2.153549171654192, 4.17123492752558), (1.7771847482106296, 2.7162852010717984, 9.477530608540238), (0.8331836551317895, 0.9292369983980786, 9.275617953415988), (6.584734077126604, 1.292638826197533, 5.633294811409692), (8.97871466865192, 2.6079923110015777, 1.2361435760068784), (7.42331290490937, 2.8772071962231105, 6.330520896053887), (2.58771162966044, 3.365592586137268, 8.256895621810907), (7.516588618032328, 4.948722510074866, 2.941189515686169), (5.74022874810322, 6.299168207206918, 6.238297763867275), (2.9470734122609743, 4.544160338627622, 1.5876051217300091), (7.791436343664623, 1.2918313925225533, 1.617262440013868)),
    ((0.07217533551424404, 1.1310930415155696, 8.98015872468741), (2.717326458193358, 4.5678163855139875, 0.7362420969840278), (2.442312617629482, 9.08155442076369, 9.33453741883902), (2.7329558959262625, 5.461810390533976, 4.828575614763585), (4.490564591886919, 3.603799153396313, 2.4143510678448035), (6.17258792997392, 5.9813437485247505, 1.8242759906350259), (1.5643292976376721, 1.0364412641547327, 6.136638118423013), (3.650596255017579, 4.325252091465383, 1.9099058618149467), (5.571498302851609, 9.358386875227572, 0.26667564791941545), (4.589842098411957, 2.5378391148447865, 4.205589687770221), (5.193884141181762, 0.5587416562110414, 1.1205517759533434), (6.4744378066193224, 5.188414628287132, 6.879531629709658), (3.6016328150115537, 2.371582424111617, 2.2949340457184175), (9.017514163385124, 3.702623628919576, 6.2992822179525545), (9.297787861555927, 7.956744736667577, 3.4322552910037976), (4.8612486412353775, 2.560982306415335, 8.97089962431224), (7.260951967897812, 1.6076494100358762, 6.716279597983837), (3.341733397793354, 8.151173022140831, 8.362462884178012), (3.6955875485939527, 7.747489139167447, 8.812408939354917), (8.629580334215465, 2.104845297228226, 3.4766216763768334), (3.7134869963018637, 8.60531317419552, 6.909103149341814), (4.468665052982943, 6.165302453521142, 0.9285287470545334), (8.722046737856594, 4.244724330453428, 7.614587534105804), (0.8636188220194463, 3.7883591634085043, 8.906492933132785), (3.2932988467305533, 9.503663539398184, 2.5843972351396016), (3.4560990449355145, 0.6604778392832633, 3.8196290510257214), (5.9818760900174315, 4.314492363236585, 4.983638898756125), (4.196955698182046, 3.147617232158443, 7.845231602351981), (6.096349423225096, 2.511531964389395, 3.792491705871445), (2.009371200065788, 8.82956608804436, 8.880277730754887), (3.72378043230177, 2.203815539564491, 3.5709168529823754), (8.5685325031545, 7.08850437987092, 0.9860471366042212)),
    ((8.106416488976752, 9.763080395993784, 2.1923465121285), (2.8002854171667693, 3.8976737180432286, 4.098674127758123), (1.2148357319983993, 1.406843451878813, 8.953504841488765), (5.339949028709247, 5.312268508178728, 6.060797109516043), (5.94833216713451, 0.001503994984581869, 3.17372824626145), (8.29957525395771, 5.161680897936013, 9.919900748709061), (9.973801871641575, 5.613237144806651, 3.538267830860302), (9.53983357488826, 0.10601641119235783, 0.6751264084809538), (2.232766037651115, 9.940684983139171, 8.787558212299588), (2.301201610894823, 1.235866134310234, 3.4068441468293154), (8.508149988812981, 6.371906024414107, 4.131060158974375), (6.548408191551394, 1.199789883823703, 6.942422665082625), (2.117750744645516, 0.592105227173938, 7.72312295923975), (0.7524873514639174, 4.467922270585763, 0.8927769266704955), (8.594017830120551, 3.3840177574175065, 7.061383867712259), (0.10139503025666907, 1.8592318676895192, 2.3892851591279163), (8.219741713049173, 7.026388879139628, 9.252880267953799), (0.5971758731809829, 1.2361942485796318, 7.038210885431284), (5.75713769810776, 6.782071067629797, 1.8497257531981626), (8.23320426641946, 5.074690589010179, 0.42683239556524866), (3.8576536385590776, 3.439154717633912, 5.70762951850578), (5.765895726186766, 7.113032082597246, 6.1392976564730875), (6.129671346572811, 1.6047860390261237, 9.81734868915513), (8.845538603205549, 8.175698136584513, 5.927088225590987), (8.56243122696135, 1.1929546820168901, 6.782128967769129), (8.960937760916215, 4.167662981031489, 6.68925355370267), (8.21291683584602, 1.8379204795198978, 2.2900877186986768), (4.474155952983983, 3.8748157259779505, 4.851542818361625), (7.863263434991205, 0.6852749522703305, 6.684408383397535), (6.691217545499729, 6.390655471602042, 0.821290069807018), (7.517391776238997, 5.691425377537388, 8.112983504817066), (5.829493077544039, 5.483332723631906, 2.603924764675977)),
    ((3.5581737402660196, 1.0952925606327724, 4.384279332241563), (6.8471674872333965, 8.088854250108316, 8.349807096945344), (3.861472774479032, 5.42490210673357, 9.836230931294745), (7.616364939401931, 3.5328002859937326, 8.714076393592663), (8.1581389362733, 4.336840960778221, 0.8334698380516725), (0.6834377985198825, 5.880027301088648, 8.690064417445615), (7.063677094684422, 2.39918862139054, 2.9715107905730265), (1.7891266364532754, 7.949134901057791, 6.452245811237393), (4.713556591286393, 4.576400504897843, 8.17071355768649), (2.360042807159126, 3.8725765994622865, 1.2159163495652159), (4.542764907103827, 8.613552913295464, 4.041282235777999), (7.583481929821431, 0.9395997696476066, 8.08430124910678), (9.798731125243684, 3.2177679928831218, 2.868734381178335), (8.373810774606186, 5.314706587361377, 4.257063863261559), (7.945806883014999, 1.379729346366192, 6.595480868545605), (8.443200416476747, 9.38856151681659, 2.472735905494672), (6.758491541705956, 9.18135617619827, 1.6121465254926515), (6.3634521020716, 0.2912161048346795, 0.9909996454262793), (7.154732010206449, 7.7157322134343165, 6.471082413707188), (6.84599240909052, 3.8499554167550185, 6.825471291371045), (6.278465827264094, 8.964231746444568, 1.8897617180794157), (0.2620663325894501, 8.907248862345082, 9.481974820771798), (3.8606972094079293, 2.3146202924603134, 9.783311529180963), (1.3358749422972815, 5.717843290360996, 0.457601923297013), (8.470929525256135, 9.312037733589358, 0.6272283963343461), (9.33521641109085, 3.2740953874138548, 9.746023626431446), (2.288003104428152, 7.963955038910156, 8.37031955635404), (2.2709975324561005, 9.908971617202685, 7.931935289267092), (4.826226654747757, 2.473050312578715, 1.7938609663065996), (4.728979201543305, 1.1026140109319393, 3.8130696650355267), (1.211766356678956, 0.005714720022939046, 5.225524808149595), (0.22016033519355216, 5.895674801957551, 4.7723302676875505)),
    ((8.727574634185357, 8.627815479406621, 7.843829197507439), (2.9381592994749006, 8.256265975330576, 2.5440577028990474), (6.224762003027941, 3.8419662115886135, 4.378627054363225), (9.181009334742633, 2.338159334928612, 9.964952481674432), (4.430123107453953, 6.798881281271157, 8.199626588981516), (5.743620830489531, 5.148884371659351, 3.8492733969931567), (2.2826170600395725, 4.2971126954420535, 8.063684931183133), (5.393667410406268, 2.203151582515207, 7.612176295123177), (1.0514716507145572, 5.593841009238263, 4.84996556978296), (5.240766748517146, 5.1517601861522895, 9.019774183465493), (4.245805244515351, 8.225869351441107, 3.63673367442337), (0.6799652250464472, 0.28098576086117766, 8.316014631654202), (9.198100993120791, 6.927673312092205, 1.5712551709564881), (1.419494923550595, 7.416251033336811, 0.7088765254055973), (3.0630153760823076, 6.215564480855411, 1.7828961214354055), (6.116510342702579, 8.333458977615296, 1.055939028293349), (2.5172991033619843, 1.7926137070288428, 7.323020454334469), (4.659635517209072, 6.549244700585961, 2.4673901500379225), (8.528830892852719, 4.785671389738982, 9.8016024385712), (1.3408623970779188, 9.101324721460896, 3.538054463219199), (0.5510389542348937, 9.840127246736884, 0.4692981413206798), (8.190134965628813, 5.663944102028151, 4.923656827948738), (7.883035491843681, 3.0310563171587255, 2.503676350029579), (6.682571803059982, 4.207884911800433, 2.5701069510814345), (1.37995889466776, 8.090591743855013, 3.661187963768157), (5.087398692325568, 9.692815497295719, 4.401399960627266), (7.040670703059052, 4.471602170989307, 2.6832809927599763), (2.138002637274238, 0.4813911482534883, 5.698946086082631), (6.700540258650638, 8.952121087918396, 6.430628183729125), (6.567109258089405, 2.487271108552951, 5.52736379385466), (1.7832233562076905, 8.308572685293408, 3.675118405552956), (5.893721928182739, 1.6064415369752871, 4.337015121636096)),
    ((9.977493803609988, 4.5566870465489595, 7.855220855038568), (5.7809358552347785, 4.629840872793642, 3.847773561732893), (0.7014264105260859, 4.217849918877393, 1.6469556225708104), (1.9311620605521962, 9.65673871605673, 5.0883231013267185), (3.639378931105963, 3.062678720258859, 8.559459726974257), (5.599083241947883, 5.689883578713028, 0.3758994148816597), (4.870629727200958, 6.438333357883241, 2.1590137802159726), (0.743192813779836, 8.04519907622701, 4.223837459860799), (7.7400264147071205, 6.708100504249144, 0.12393994039224032), (4.054913168800161, 1.0427197726405502, 9.696603844201084), (2.4242011599595314, 0.8088435784285763, 0.42817775088326737), (2.148078136197511, 0.9875788889993464, 1.657991270541952), (8.57080318648859, 7.132573887127612, 3.124175570490386), (6.254344422255258, 0.04871096137175068, 0.9567327772703016), (5.524060147480752, 4.317449436595588, 1.9056409490653414), (4.208479300490351, 1.0977166857611875, 0.8031109128860414), (2.8388366796510156, 2.505983354327136, 9.717210024646075), (0.7030296926038415, 3.28850086554324, 4.75908395274661), (9.550798468931754, 2.719523699317082, 6.238275091224166), (2.1496371326388832, 2.0529632522918115, 9.774436559148285), (1.4690495307973872, 6.080277879483322, 0.046337383939615284), (6.37675006066517, 7.516635540272944, 6.1165130891621615), (7.999790319294737, 4.016194640676112, 6.575816053558339), (1.9053555340856954, 9.824253933151674, 2.4400403247764513), (2.2530941931775206, 4.945193630179583, 7.659347084349763), (1.9102919021017084, 6.60919685686138, 1.2339653022973163), (3.689965303585958, 2.407862731456656, 5.119316472008188), (4.231046873633884, 2.4160468700264737, 4.914478801593542), (4.340004636968635, 2.332913875023589, 0.9074402484443245), (9.359461283697929, 9.290851533790404, 9.720315936411136), (1.171163220134036, 7.963309680337697, 8.770010609283263), (4.004155322260842, 4.8887211747351245, 6.7335963971237796)),
    ((1.3265864160213259, 3.7903739745935674, 2.3184587215643693), (3.1850439232861607, 8.792657330020246, 2.2508318917712233), (5.711056269083526, 4.031534217211517, 1.056337164721094), (7.06106630849677, 2.232320928381996, 0.17331316762925764), (5.236254425576998, 4.079839602294331, 5.94014607318991), (8.246876546297635, 1.656792716181279, 9.044862125749317), (3.090569413945665, 7.177576336939352, 2.541826553845584), (2.3932664869723275, 5.863622757700205, 6.448793136608462), (7.422851304290957, 2.9260029458521917, 2.8892356421848673), (0.8754738450237531, 8.109759389650863, 1.3139961385812249), (7.058688111292507, 8.339180737283074, 0.9819372087849954), (6.643782395351767, 9.536899359322428, 6.356482634064113), (0.9679684253666287, 7.580335551284803, 1.7793725108717795), (9.666255679325278, 4.037532584925768, 8.149917697231434), (7.084542471054701, 2.012873457439764, 3.9072860429422676), (9.920424430933254, 0.2161226098262492, 1.4318465912550349), (0.39241996700773885, 0.7315000861534549, 7.197863547655059), (5.1672234533828245, 1.9255407124464097, 2.752983637757901), (3.6380146711028827, 4.143495316257496, 9.839024913366663), (1.5676958117237494, 0.7222032245157639, 7.188129461847264), (0.7905186169240475, 1.8660276220055905, 7.833336196375922), (0.6141542410535494, 5.9431616081872916, 2.921951869044653), (7.082396846820416, 5.588437033152928, 6.160834436817292), (7.374062307492146, 4.59736909100595, 9.243617653050997), (3.6417292591583528, 4.401032486297409, 4.355529897289413), (8.371075042964343, 7.314424970850959, 8.656087319592782), (6.986959546467343, 8.564752620721366, 6.320937975471538), (4.94969745722991, 9.533146360725151, 3.1035337321581844), (8.980004199412733, 0.7288860655877549, 7.6945583949397065), (3.918528807197813, 8.154479703879186, 7.224632944767304), (3.373305193091869, 3.5347225190035125, 6.027616400290223), (2.4931935167588315, 8.226251821468267, 0.6460830591987421)),
    ((8.805205852578382, 5.206820117196676, 3.755817497388414), (1.884487081543611, 3.6073353613116366, 5.457958453357671), (8.965727218329572, 0.09827577369057039, 1.5300480196528332), (6.939941915760369, 8.754652373038306, 9.61044552888524), (4.334698386781042, 2.0960112423563295, 5.754602266251352), (9.197579140083503, 2.7665611489347097, 1.4470287149606331), (8.88514684809525, 0.801212941343421, 2.8383342641675444), (0.5601317047874099, 6.584005652230948, 1.810023958939967), (6.9221260330459415, 0.26243966030387034, 9.10690695813425), (1.24606127035922, 5.602902623402634, 8.680823098483351), (8.923768987147444, 2.142332414577175, 3.7597786867155856), (3.6745235621179195, 5.047061926355846, 4.0604590541516306), (7.658761361060843, 9.183414453902182, 6.0033284925518355), (8.701791004080029, 7.235105063914547, 9.687632915591069), (0.012852190718217749, 0.856715796229055, 9.111976743358092), (1.9594302883735149, 3.1203579397049417, 6.551966447140646), (8.439568825794305, 4.549976489865189, 0.7571427153739996), (0.5569674895480581, 4.147972606494854, 5.126105175592038), (7.5496184931659736, 3.057620845654779, 5.541498316233636), (2.580491211582745, 6.228613889610055, 6.341451227378046), (8.229344996263418, 3.443714192394883, 9.09597312223155), (8.46171419791816, 0.28189008064609, 5.689727273416781), (9.102705615194553, 6.271202169759765, 5.833586686998621), (6.940137472375364, 8.303312496921533, 2.5287082681516404), (7.668272671744099, 1.5909073419160014, 9.000751392521087), (2.3894901264015287, 1.3560791273040196, 9.59900558451945), (2.659597067734718, 1.2613612903763949, 1.6820695804517982), (8.2344705462326, 2.2270052413716543, 9.121378925999945), (1.3599227075163878, 2.7499175606460713, 5.8411143487888175), (4.144394732295998, 0.6379444170784454, 3.7353940027829835), (2.4913361276047885, 3.175423217439979, 3.923898538353827), (4.396616113795097, 5.537770744156988, 6.873463858307414)),
    ((6.269990775595105, 3.9547358809721347, 6.592174126003764), (9.798690615743157, 0.06574531749882206, 2.6895618967245993), (8.230706500790808, 2.9367694428004345, 4.543355783406884), (1.411146633793029, 5.132056380110753, 3.0832295669409024), (8.898699736144117, 3.316064846663619, 7.29161079668407), (2.2732660549267436, 0.8942634450511799, 4.241293997565765), (1.0828313433535686, 1.849885389008793, 7.5700777417726375), (8.870429811809592, 3.456366620360968, 1.2054609399128446), (0.02360933508824714, 0.1650723698321943, 3.455684369967462), (9.886990852139729, 2.256303476655943, 7.347802029762091), (5.92080056421336, 0.9081090737045805, 0.6286456331289403), (4.171932540974423, 7.217581313891581, 9.951478544273364), (2.390245454052536, 9.417030370709764, 1.2673084259396117), (0.8647812162741919, 9.408810226950301, 4.991730671037644), (3.9895622360571767, 7.0202222993806584, 5.8519832303152475), (3.877404449900558, 8.040533163201511, 5.288789666436015), (2.8104310945453115, 9.384636821213492, 5.57240296126278), (6.152326636260107, 1.0407413845395252, 2.3628102098352057), (0.28417783868183166, 2.459292448255707, 7.704208322747082), (8.403108627903897, 9.170811979015843, 6.917426131340669), (2.9646199280325822, 1.0189639209676105, 1.9404763634073985), (2.8164473643532393, 9.088684197061541, 3.1806452637585005), (1.3949818446403106, 8.201722005326564, 8.240456133115106), (2.2683752905863184, 2.703337209539416, 7.328332015386136), (7.029723108823794, 8.064722641083998, 9.183443781794068), (7.641252805165578, 8.518957454034242, 0.4602026842071305), (3.5612058384798786, 6.8932152733994165, 5.799793639566689), (5.757970756690154, 0.5828532321758617, 7.018930402689443), (0.8578393234331827, 7.91560269636568, 9.363255449771792), (7.6951976050958235, 7.4271751443054566, 7.496266505242367), (4.309706188798808, 3.981774425700426, 9.214862616707567), (7.116105955457799, 5.473386233416219, 5.795661427850884)),
    ((9.134415295420386, 6.525291387814413, 1.072131278955989), (6.297779689228893, 3.640313373044688, 7.510300977202635), (6.560075686275263, 6.589072578922421, 5.682326574743975), (9.482184342875208, 7.358810641866675, 2.9951564928325833), (5.486528037633435, 8.73183702577164, 1.8337785855500621), (6.44937692355974, 7.488477215902579, 2.2134871045459157), (0.7239654471904189, 2.9370457770266736, 1.818179485396314), (8.854122163351585, 5.913701875222907, 1.7115972885278408), (8.800072427701558, 5.757299923742181, 2.1446873547884246), (4.565019929145603, 5.2870785592410705, 7.268018078934272), (4.579967323226105, 1.9352967337232319, 1.9330743194021638), (5.782948571029384, 3.889751708566446, 7.348549240790973), (7.400511100643325, 5.411435160818312, 8.34552099576707), (2.156401503076885, 6.432397333062792, 8.858396257258592), (3.8102445994561664, 1.534011000513117, 9.00899264857996), (3.343870897867535, 3.0161889404665887, 7.952061420616488), (5.04498842597345, 4.700827258204809, 2.8487427112643484), (6.0889164066516965, 0.03950822704847812, 1.3494788793131296), (9.919968203753717, 7.385881971922201, 7.336607554020006), (5.115476820098462, 5.880041692522584, 1.4008305604561089), (3.428851161873503, 7.1817195085045995, 7.527488252530491), (5.6221641998747085, 8.430099015406675, 7.89920101129132), (8.424129348314011, 4.906245801210654, 4.889621546829405), (2.280658029148378, 8.70008945432584, 1.156751525954649), (4.322768753618905, 4.200922081354141, 0.5994820781801735), (2.402395345115912, 9.884588407563182, 8.007207665089076), (6.940737840379674, 1.9736228967823333, 5.074178481533721), (9.535683997898293, 3.8224101661724905, 8.422914350832993), (1.4294058634766516, 8.863641521031047, 0.37820330904697497), (7.815706408544983, 9.532452955733028, 6.27949019255865), (3.6660372958876697, 1.8703437648009158, 1.614839070885865), (6.405518927138347, 9.697007320141648, 6.522679757871959)),
    ((8.642217639647349, 6.196298109853226, 0.188782324261193), (7.7770204624093795, 8.322413402186744, 3.470770579634647), (7.124038603361211, 3.748312409923773, 7.093929841142258), (8.820650186055873, 1.5997245654818049, 3.0085134051915063), (0.5483722806913816, 2.8178408616073822, 5.706018852013905), (5.1145873684524705, 6.80917061203333, 2.3033398627494464), (4.332677738161107, 8.263830982335683, 3.5711577266240724), (1.631230909837157, 7.005687861380988, 8.982360842021608), (9.800603433305774, 9.09617022304285, 6.981754300441494), (3.6868455939173153, 6.285683090438506, 0.1683906251137346), (6.6042656708297365, 7.886043152067139, 1.9137166040699038), (8.054357602275001, 4.421064128361365, 1.650723125244794), (4.060021152094997, 2.6906350910405807, 7.756959413215439), (1.2614505813936683, 6.275776758360834, 2.451351824590952), (0.33793623357379343, 2.0867778043086616, 0.48281356152430677), (6.46049900335263, 0.8064155136819773, 7.686960606401843), (3.0403818031465137, 1.7642469095491764, 2.368046326298722), (1.5103867216815103, 0.02656423887319681, 9.754401363680183), (5.277923028008172, 6.030917580545163, 3.864086477696601), (5.175479862537829, 5.076934488986136, 2.47992503328069), (0.570651533584613, 1.3971647846821322, 6.348787842795111), (7.922003320586373, 7.646254359279085, 7.273730883402871), (6.722479731321696, 8.033943849026489, 7.165744708396532), (8.882760513096253, 1.8181072427106248, 7.174677568583125), (2.320812123275947, 3.632287872155687, 9.860865316055348), (9.96237601114013, 8.35653031171651, 4.428389060100379), (1.9410072070404527, 7.008457701582019, 4.188786728567354), (0.4050859939535656, 1.275878087401675, 0.9658562054504438), (0.9562387637091196, 1.6841865201833695, 0.6933058045683815), (9.523603198135103, 0.6311505595011035, 7.28888787237274), (3.332278709899681, 1.1859705224354389, 9.201595342335565), (7.572785089227763, 9.688927358855743, 1.4440756800728438)),
    ((0.803246043130682, 8.678921249935136, 0.6171211079038608), (7.421846206773682, 9.96606133280624, 3.7122102385829727), (2.9960069148711552, 4.101250790377265, 5.527680912361768), (3.113910006374719, 1.1659120171673287, 8.270138641570512), (2.330834081965114, 3.0613495115926073, 4.113642249507978), (0.8515123045011519, 0.7582515492948805, 7.350660476333456), (5.916011609297136, 0.1883266234856551, 5.725726432390127), (1.6939446343212294, 7.6325030134540475, 6.372521765035174), (8.796516792476645, 8.18502806201765, 7.888118436679303), (9.251758735271768, 6.679049304994887, 8.163203963498072), (5.248959689839367, 4.89989557860301, 4.211160124734885), (3.808626641819748, 3.1532933780665493, 2.442643510630754), (0.926914591794924, 9.757276219806824, 9.726358807611245), (1.6616503301226448, 5.035823467031198, 6.339789405364703), (6.10445524448585, 1.4436073569798802, 8.742516303211618), (2.6090600494477667, 5.530270722999231, 4.810414493258989), (8.017439725302697, 9.658818044205368, 4.160941917930229), (7.078991192950199, 7.332586264141183, 4.726405420841724), (7.57641746285617, 6.349557291591459, 4.7856215235130275), (1.0598633928889245, 4.048872457978515, 1.9001534781300289), (6.214813908717107, 4.548061767639419, 2.882007641256066), (3.9139685629743126, 8.633688852108934, 5.229943376613074), (7.334110403852662, 4.454548086495862, 5.196191307509624), (4.790980737902326, 6.115058813647119, 9.270422685405123), (8.185791887597308, 8.189375909640027, 7.549102432948576), (8.903218159390985, 8.205839562082483, 7.713887269365881), (9.440851665215815, 3.601670947374541, 6.48124509023731), (2.599402239588878, 9.377751910999875, 1.2988807799763369), (3.143693902273088, 1.1971122980816395, 6.504367795170936), (8.42000101928822, 2.4689811356631908, 8.21824793682127), (6.468619521823637, 7.828147389335619, 8.75189764096186), (4.974054043584408, 3.1585661510147514, 3.4794532707038783)),
    ((2.3886701993910853, 6.388438042448134, 2.9102788254295566), (9.531749961993892, 8.217505194453746, 7.233521577292297), (4.048381227028317, 3.654340747304623, 1.5954556226449557), (3.7924318619599684, 5.8775223591263455, 5.807219580351153), (1.3604460026216136, 0.8108513126490724, 1.4214554013252245), (6.405289886634201, 7.8512680044074905, 1.4225330319779117), (0.2914722327865982, 7.988686562520014, 6.854162574064173), (8.365933560708045, 5.5864550735405505, 5.27092689567737), (1.1524217608684406, 0.4005868812801838, 6.3169929171233585), (2.412240422732838, 6.5336862335731105, 9.246858908306674), (0.678997193278188, 3.016886339112541, 6.199417505407419), (6.739793359625943, 9.172889110784979, 4.59266536158657), (1.34788850580851, 7.4567420548683305, 4.2768260425573645), (3.303686749182515, 6.369844046096896, 5.244880918174088), (0.9055911731104005, 6.523753122108021, 1.5316887474619723), (9.698433498615284, 5.197206939709222, 1.054592775063613), (7.702599299867292, 8.719242270997603, 8.743913291639346), (6.642634938068818, 6.740204120834708, 0.6721977027010395), (3.1968249589563658, 7.227132029318141, 3.8822376141345805), (1.171707195212518, 0.2962629278430484, 7.838017826894838), (1.5133243859392365, 2.6506639657420483, 2.582657541389911), (5.5000660297053985, 1.4876336579112037, 5.443455489422629), (8.272143810551643, 0.9311217798272386, 2.5566583402989185), (1.964734809615134, 1.3777174352297639, 4.671722123854777), (5.535020581506328, 0.4558701750801386, 9.41121931481009), (2.5900759771055473, 2.289456625813439, 5.458324566030965), (8.237331902499607, 2.558995132391196, 5.207963770941734), (3.8759106275684885, 1.1240938334304151, 6.179341740535909), (6.011136288788796, 9.170283047854511, 6.079328306127301), (0.7167206382619895, 0.8067838551172724, 5.7484705271402605), (1.718545197138136, 2.7241312599214784, 0.5592698878377012), (1.4050756314062973, 8.96360549014385, 2.6677230691850373)),
    ((1.1402549925570116, 9.971978151673135, 1.3570350932787956), (2.1389901427426636, 2.1104118476753833, 9.645307671280005), (0.625458380057835, 0.8270695896578195, 1.4985525333075111), (3.0673077265636595, 8.638105130117092, 2.3703548231337512), (8.701649959887101, 3.9070408300384054, 3.589856922069521), (5.074089065441635, 0.8540919760476318, 4.925773747237083), (1.752411275116884, 6.839358635233505, 8.716205729828623), (8.349438912759764, 3.9142116394320006, 4.838373772819967), (5.15025553915839, 3.070558575820048, 4.231753018460398), (5.925960064028329, 5.904012188875686, 5.3768095361269275), (3.4514768137465435, 6.973071761104634, 9.435518061392719), (3.384082049222049, 5.9922807780583955, 3.3554399275197886), (4.378966938477246, 2.6408852253798756, 7.301263720571599), (9.97762077329149, 8.844756450247962, 0.9911624998391166), (9.853099833402414, 1.1966178248438253, 9.206501858260998), (4.0251329468873145, 0.05269880378702241, 8.533976792138684), (6.310787404625602, 5.595255074384568, 9.525304498911689), (4.931428173155547, 3.377532388300166, 7.720572103273621), (3.032529804339995, 4.380073036829528, 3.5945949157375088), (8.386882306595773, 7.629924929929793, 2.2344313361170407), (2.0155769357427133, 3.477514260398199, 8.745279286112062), (4.049006162214363, 7.1950262469316595, 5.195454066252658), (6.956481143537058, 3.585480002102832, 6.935763668440633), (1.2143004909213484, 9.872583104354135, 7.826376321374166), (0.6107407681990551, 6.812157640856138, 6.822008458785104), (2.3072347838799914, 7.498523114721141, 4.109557318818355), (9.35856164437332, 3.2667661587720254, 9.110385140342476), (2.2548467598475455, 9.22700219580297, 4.783312715040628), (5.455945049149693, 6.267437033319812, 8.168865267854398), (3.993844685595429, 7.4512721128614015, 8.132564147814959), (0.8895108655702577, 9.29461242597797, 0.38981745573915316), (4.75358273201728, 8.925374519388443, 3.312474256930771)),
    ((3.6874847569529257, 0.0660401692088497, 4.123274859389898), (1.3829970156510552, 1.0724060867565655, 7.247368080113903), (9.872044260142914, 3.021938576207649, 5.406486824605109), (0.9593555495136985, 3.8275274851666516, 9.547207927459956), (9.601222562568344, 3.392967972801056, 6.324709590956412), (1.5319796364963933, 3.062679529545097, 7.126743732699169), (1.2084735202451524, 5.851335809619526, 3.8523597534300524), (6.232220383675991, 8.991035564189092, 4.9519926926747555), (0.22665276916125077, 4.947420213223083, 8.25590912207398), (4.0466656814899435, 4.037232758235253, 0.286132961502491), (0.9715089576677027, 4.1166682181964624, 5.79625018399761), (7.580512295505458, 2.2024722237905614, 1.2719259466653676), (0.7623435019622105, 5.538051385989445, 3.8953441616198834), (0.1317896373584182, 9.525394317603977, 1.6381049466988928), (8.701739776735032, 5.563810345714602, 3.756024754282541), (7.6607734526407345, 2.518795804495114, 6.960320418930937), (9.662499927104452, 8.677533617133825, 0.7480072131376225), (5.491976346393905, 3.5919146996916087, 2.22694536631731), (5.647877103392461, 4.438225916367498, 8.692152598657586), (2.8481377774661443, 6.000518851092678, 8.002550259855715), (4.307711439479473, 1.2896582812153579, 2.7304861986965423), (6.539765376185902, 7.833874648864832, 8.070529685986859), (6.129014482925834, 9.99429677895262, 7.191310144656931), (8.089378582450342, 6.759352111540201, 9.040157873265068), (1.962828981645538, 9.369068197988838, 6.514734718737667), (8.15015268141249, 0.6324014240523568, 3.529103328072114), (8.622407585109658, 6.888702277181532, 4.69112767761111), (2.9906546986108964, 9.233409119997619, 5.779946102849726), (0.6476735102874276, 2.0642688881582636, 4.504929630079836), (2.3219771157977833, 4.842742419112739, 7.835298073936646), (8.365687739323882, 3.262903759197026, 1.2735852150295623), (1.0812536529088457, 2.4805045434134176, 6.347211627838791)),
    ((3.9415650645743683, 3.531340915180726, 9.152124852530527), (9.137505180254992, 4.083317988230575, 3.233744935249697), (0.21055940044144017, 1.641248068788952, 3.72035174653179), (1.58843604321118, 5.477970318998681, 3.394029441492844), (0.576356327749804, 5.139552732510625, 8.287821169981935), (3.667391451481773, 0.35082582670492246, 0.5618316890213915), (6.250291486008862, 8.852437884629312, 7.420088765488009), (7.567601105782562, 0.474043933460806, 8.03969862647104), (8.182058142248241, 9.886946836711733, 8.9091520010359), (4.354324251356249, 0.9089513121193238, 7.382430530938859), (4.919517813053628, 2.0424311017660224, 3.721710182294636), (0.1354471552753933, 7.698069742776873, 3.739194434670572), (1.508523276636402, 0.43925419538626165, 2.6287259453066225), (2.9452355471972957, 1.975700083891806, 7.989992607695839), (4.0219083406150595, 5.960226417727078, 5.914622711353025), (2.9696438073420675, 8.639675663589239, 7.7459532308694), (3.0631547920970736, 6.54248204714626, 3.551060207146027), (9.204234773519806, 3.027035693351272, 6.904181750247719), (8.925610368244932, 7.664107179019329, 6.5254140083687275), (5.029638898575004, 2.32862279745774, 3.6347816275339673), (5.942025250651871, 8.212644309074971, 0.624058458672897), (4.569878988458752, 6.491116138662608, 8.098463091726323), (2.6961526860966623, 5.466216050700462, 9.613431426941334), (0.12496485649828637, 6.879010260342273, 5.103693763947086), (5.939405424339418, 0.36990569424281916, 0.22985622593195587), (0.38941199759941814, 0.9392931844159158, 9.618501693352687), (0.48339797243360016, 8.291289280303197, 9.353941341963516), (0.3700526161670614, 1.4678148875703023, 0.3911510362354298), (5.329667512084795, 0.45539217334750415, 9.728878535774081), (7.6286119392132425, 2.290371280990499, 4.276051243638923), (4.889481093342587, 3.123872200768112, 1.4673977019058182), (5.105140785584434, 5.808007734763226, 7.781954136673761)),
    ((4.885887841884782, 9.58452323045217, 4.038849803628873), (0.6191365079961997, 2.796239139776091, 0.030395540420438127), (2.4488456382774624, 9.835658592133715, 6.210078968851034), (6.510997247324246, 0.6538533402781677, 5.110305709650086), (9.735284578167299, 1.6965517891051474, 1.1206305314553633), (6.205682834382599, 4.4009595865874305, 9.60031011942202), (8.005197645744985, 3.3540822845792695, 2.131575984558091), (1.3970990772677616, 7.484723618794662, 3.9556163911900653), (6.28483239394768, 1.684590328077722, 8.719655915280383), (6.829188240309236, 0.9771623284828668, 8.603538879122004), (2.2669983379862355, 0.26885621064440146, 3.458674483885039), (8.237708693106132, 0.11363292364556132, 6.697783419834627), (8.09899591825265, 0.932188969442731, 7.778653330970204), (8.472221236277921, 7.008712786720458, 3.026644062610775), (2.4026666801455256, 9.197303175438824, 4.659498260550271), (0.68478363626581, 7.181785377191493, 3.1896760804077315), (1.5933852376890922, 9.192162248185742, 8.899125174580554), (4.244566104823853, 3.411969368312354, 4.24787335077892), (4.015045230686902, 0.708448232301, 5.429565477278613), (8.458763451658687, 4.195104793887495, 0.6515652928779692), (7.827544319947415, 0.15096692511333276, 8.716617171138028), (8.59777753028567, 5.7912542641518385, 9.761716463316674), (9.62233983741275, 8.261740480502818, 4.811037504486872), (2.9190535658356023, 7.965650457670602, 0.24285460616874532), (0.7473967595587239, 8.465518858305357, 0.023828579490563495), (2.0287767821692393, 5.329504661221486, 6.590013349779013), (4.022351002317474, 3.9448711618435084, 5.638296883041507), (6.299731629364711, 4.767576059200268, 9.591794109898206), (6.879659927383736, 3.430052810546255, 8.816899477597888), (5.372263013759035, 4.57142749557888, 4.977031660296525), (1.809940718093862, 2.0393392456861137, 0.060833710531928986), (5.226440062057693, 2.8654096484691816, 5.740604889781532)),
    ((6.852087871089113, 9.108313960921192, 2.2183177404100918), (9.274675123996346, 3.947779924816106, 9.661035574351605), (9.40940922106254, 7.890818818373844, 5.57590597258459), (8.676842134678438, 6.375979228542793, 4.535890869365822), (4.351429148397634, 5.543539456620708, 0.10839394680602465), (6.1969234483257685, 8.303708653086284, 7.966084647675318), (6.63124276418578, 6.893946409962681, 2.5347149415231085), (3.2378339530463163, 8.725363100734624, 5.293426810331479), (6.4689630846873145, 5.050539866461159, 5.7153920268115765), (1.7661648949522546, 0.31439926763757287, 1.2211255131368548), (6.133194512095691, 0.10295601755988426, 8.241960996857047), (0.5357128892345631, 1.0610337860995556, 9.89042740574616), (1.2231738600341024, 0.8667800061776387, 4.004530349634649), (8.678377422067095, 3.318506365759962, 9.586037107303332), (3.569728101802907, 3.845840564678167, 9.118506847110934), (2.2958138746341006, 8.402721247727799, 7.214290173342214), (7.912494572282495, 6.401826872375249, 6.894802738984193), (7.309900591510763, 0.4169859100943718, 1.1373442591044647), (8.984711429819544, 2.619239118070614, 2.3947397779361057), (0.5030538588563749, 2.406821221338864, 8.301613486538427), (9.134171892749489, 1.977841967602113, 9.301467547623801), (5.099001355137273, 0.02716435195165734, 9.169719107163592), (3.869595193420854, 0.4886389111863354, 2.839388415459436), (2.4779712662459596, 8.81702135294195, 4.62457784698867), (1.84981704135171, 8.306241785588435, 8.14965557941645), (0.4274388816415686, 2.6608053191280168, 6.7016514385682315), (0.13148173283956455, 0.09722683045968794, 7.066949969746177), (6.221492897036317, 9.863806632329888, 1.1621597992720567), (9.567468566033835, 3.3169277329001012, 7.342785711385828), (1.3296258487565515, 6.435993079850132, 7.286867042419778), (0.08413492044841209, 1.4650191717052374, 3.281551675454044), (2.8202569784429956, 8.907262663211386, 6.076954250389491)),
    ((9.758402834545416, 2.8587786978921126, 1.407142117351673), (7.737051824767653, 9.804951591629335, 6.899803723625424), (2.0723068287419686, 1.3823954917068437, 3.560562186565183), (8.985767793297367, 6.49413448852984, 9.761689148022526), (0.3012740662682589, 7.468934243664563, 3.0628199391752475), (4.343131850253615, 7.752024775066912, 5.348308537308446), (8.63420113534771, 8.185313085335652, 8.398183522335241), (4.657640069777092, 7.507086707340971, 1.9113884275888748), (6.9768839051632785, 9.584660777276946, 6.303379852402138), (5.600805352008086, 5.0985144931659985, 4.47369711922212), (4.314682996153195, 0.3594026397580552, 7.542392034091864), (4.893554430675666, 0.2785042977786789, 4.882062251951861), (0.547756537152454, 1.1280590806855118, 3.3301993066074944), (6.864429490429018, 9.330681747684231, 4.258599745568916), (9.233637083130384, 2.6639464091302747, 7.37389798889068), (7.800347549365374, 3.8270479693448136, 3.5842898326997386), (6.465940796965095, 6.260566329084947, 8.934116255405913), (3.701049049855331, 1.22716459512763, 9.4002631640118), (4.693268633528268, 7.846437084023616, 4.196030407100977), (4.891949942049267, 6.534956133995617, 5.4883474540203085), (8.673878927263264, 8.688741051083632, 4.608968506871936), (3.3765762915422615, 7.589035492753462, 8.658282816096335), (1.2953328220402793, 4.247897819153074, 7.686479958029047), (8.985645237358991, 7.361325000517044, 6.674609832338145), (4.78160361081242, 2.167029367430003, 3.418518533922996), (4.903669364673205, 1.4889897098918892, 4.840183990624797), (2.656491220616213, 7.200767821073998, 4.013348377411967), (8.907411599010095, 9.485423973791407, 2.03671249895496), (3.5650683202522737, 2.6189074662415948, 6.592455214598234), (7.2150846216843165, 0.49129076083658796, 9.610042075683157), (8.677118281005477, 9.240488213137283, 4.197813436441008), (0.07237846193325459, 8.135939173913997, 7.141216286164043)),
    ((1.052079384156711, 8.077115754696969, 3.91397464098406), (9.403674392801499, 2.8677887800087767, 8.403220196486753), (8.333588598818523, 0.4682482665606058, 6.9738117131034), (2.786979345175987, 9.75203822428709, 0.5915259878042034), (3.539768851225392, 8.122053412787528, 9.793650329886248), (3.3118468483702603, 3.7751738244468758, 6.35048421949914), (6.792512518363573, 2.7770008664982937, 2.9887891745885184), (8.234362709730162, 5.271904998597793, 2.8871049474343224), (6.59060015696239, 8.88792157416218, 7.651023182793994), (4.073769563544662, 8.447440243578754, 0.8992646537457216), (1.8164288811326745, 6.2337074399744985, 6.313241966027222), (7.521017962074752, 6.699373988966454, 8.122095071405678), (6.210780739812179, 4.746574258964495, 8.221860719290586), (0.8875601301411451, 9.570253544522895, 5.247287927737778), (4.3570065324357, 0.4338350928852941, 4.882615039720363), (7.769187020022381, 1.8943647965430166, 4.377654487577849), (7.8753121749391095, 3.6771025100101684, 5.631696227749497), (4.089571857562024, 4.033952096217503, 7.762884013411919), (0.3242240554869913, 2.1118523525646515, 0.2951485125143538), (3.144654626000689, 4.703929126295794, 8.236617714307794), (7.537452401168001, 7.048601319200813, 5.9197555951761505), (8.115884192605805, 2.546368231962547, 7.856094563363724), (1.6703387195759634, 3.944602537917532, 5.5690513900720156), (9.999039297720465, 1.0815269092819568, 1.9495577736663128), (7.940593116112664, 8.003902891957178, 5.202835768576363), (9.31731902268396, 8.010674739792197, 8.668827305749513), (8.205228056467668, 5.782202921688469, 3.3537540866372284), (4.165976009726073, 2.5223155366032444, 0.5555477660397645), (5.913132407724375, 6.14409201168629, 8.267577432000689), (5.39394974741715, 9.075927488472045, 4.189534942151071), (0.5690985502158663, 0.1578582468883183, 5.3656635618187), (4.157914876358822, 6.8728835343691035, 9.584422489446334)),
    ((7.967195296393498, 8.295442003801249, 0.5520303581062291), (3.8859392824481964, 0.27880109578231727, 7.169422641710104), (2.3189225376857827, 8.859401047083093, 6.108978975196768), (1.6659311291158774, 5.3869518079507746, 4.534255736362162), (2.096546882960577, 1.0838561744026043, 4.980795903179416), (1.2251072569738375, 0.38610779197029266, 2.628634949048212), (7.277699764273825, 1.223076664843028, 6.335811759608989), (5.5109068047764795, 7.758524845293415, 2.3577898517613516), (3.1330675138269317, 2.282331833844303, 5.7909400657598775), (8.226543079005296, 0.3540109029624028, 4.007247937919763), (0.7525251422653145, 7.324512240445219, 8.7967606497889), (7.524411056143685, 6.13016090226108, 7.908501802003459), (5.792261100888848, 0.8066627382376412, 0.4147971122098726), (5.045565785893911, 7.568768383451352, 5.324841274698667), (7.828040361857678, 6.114474867459246, 7.048756543513011), (8.656721884667611, 4.671199495181062, 3.3831369030606573), (9.634150303907212, 3.0944809083933777, 9.368016148829922), (6.817311347496097, 2.081843006129831, 4.862935947884209), (2.9227579638747017, 9.748068169423261, 6.164509992756567), (2.557757350563369, 5.490378722611907, 5.532000389021963), (7.732485944415296, 7.7904821262365065, 6.333853805389654), (4.285510246234971, 7.467810441475925, 2.249807348374272), (6.068657723821923, 4.730241090199786, 2.3352008352063125), (3.5157947346381757, 7.839079268034954, 7.242492476868899), (5.5060528239982425, 5.275349965065631, 9.7336046887211), (4.064889125259205, 1.8128143165748722, 4.041803520889406), (9.614980394188912, 7.326167481321448, 4.835630103796929), (0.7346604102434606, 0.782997243298359, 5.1293489953342775), (9.425542675735821, 7.40488111142255, 5.708639555094828), (6.378370605074094, 9.023251918064886, 1.5824028950785207), (6.111848505297422, 4.438677968182516, 2.4792553788757035), (1.0984084314393272, 2.08049865681879, 7.420081864461205)),
    ((2.8586179148815374, 5.174403481687936, 2.38413897704983), (8.936905115653392, 1.3675166671596661, 2.8364041533166997), (1.7884134773919136, 0.7961762513220827, 8.470913547095618), (7.130991384942337, 6.789703767427487, 0.2458774711093603), (5.334633280240942, 7.260138292107726, 5.249529312785289), (1.564510990385779, 7.423136289184839, 5.70399058217453), (0.8915708518268539, 1.2804847100908168, 6.791935606118763), (2.2550252799429202, 3.398347581616965, 8.976037111062091), (8.768271690418754, 2.425239818107409, 2.2509408115348464), (8.598042114517096, 0.4424976491378141, 4.534878713490719), (2.9917401196054594, 7.38899492093922, 4.825581165586325), (0.6068495439393184, 8.94801024778738, 8.692312304473777), (9.936360540128547, 4.521774452361336, 7.022117136872044), (7.643417610351502, 7.538150460209838, 9.29353182453075), (4.251225864456995, 3.2562040347108443, 6.931612999465675), (3.5724755033007916, 3.762097789235196, 8.511059565855115), (8.559700847605718, 2.3585527503140113, 8.541075328685997), (3.4917683917932485, 4.31866960446349, 3.5892441818154452), (0.6517090113044899, 0.5472156947299123, 5.921760936026088), (7.762978888079479, 4.588275528483853, 6.027938689759962), (6.235139990896542, 2.088320693041157, 0.007661542379296948), (3.979379580823971, 5.679446041167005, 7.788689773722383), (0.29099081466784305, 1.6547782681254286, 8.79500194398019), (5.676711413623778, 7.763599655570859, 1.9787887034572194), (5.433390183242254, 4.149779323951421, 3.4809789197334995), (0.17063278055386988, 9.4935853081832, 5.229890054132218), (1.7634167504633202, 1.6193521416473133, 2.2404024468434915), (1.8940299709783226, 7.397957356907429, 3.1918521058029716), (4.8850107815995605, 9.377036666017082, 8.940678088639277), (0.7163030677362525, 3.672103652307216, 2.214655385281082), (6.419544735955669, 1.623994108815442, 1.2342780027068123), (6.897963022907856, 7.146654886384574, 1.4095242175851097)),
    ((9.596869435047243, 1.6971622119622831, 5.471559535870121), (0.3658360035251984, 5.042143640080846, 0.34557807384268835), (3.6643271198780383, 3.156869216828518, 3.956199484972327), (4.507571704282389, 8.587800492904044, 3.776916601764777), (3.8024626430667596, 1.6812544282277653, 5.850859318500834), (1.3164734644545573, 1.007956095056599, 4.823993486852824), (0.43744211502286356, 7.729783717139492, 7.9120214818271855), (3.0999223334149417, 9.63100672359299, 6.161780931908849), (8.886063576066803, 0.7185820530189779, 1.2597934022129742), (3.747654492523761, 2.6130997347814064, 2.971500018108446), (5.918291732230569, 2.724214277066641, 0.895325188147833), (9.631805120580175, 2.8470787895448737, 6.983586590078067), (3.8134221807946336, 0.477646053806714, 9.485355598164322), (8.97850940600156, 2.452370933357458, 9.801233058426899), (7.484220249734804, 8.109538877762114, 7.767317316247172), (4.51927310990905, 7.360719488969424, 9.981326321435827), (8.826147747787799, 8.165287354076867, 8.631379723593275), (2.5074609948263484, 1.7118905484125313, 6.02502509400074), (6.99220184486264, 3.7158737559490085, 2.6704218862402387), (0.3623826834672428, 9.841919335919052, 5.2744487148428405), (7.401870290499946, 8.129082092079035, 3.669339711865105), (4.263514020277094, 9.80838017177134, 5.888696809779378), (0.04318800025939318, 8.242374419167925, 5.91025983943948), (2.890015649447334, 2.097471182682331, 0.42691792632057135), (5.65738067369495, 8.01636379334142, 7.956156913847234), (1.765209704314522, 0.7640093498348599, 0.5697884644841511), (8.343467590843064, 4.367329109835698, 9.189198614795952), (9.481527303146725, 4.100959481288404, 6.5158422061774965), (8.190664020420877, 5.816073051401958, 6.546070578002114), (5.784246667526068, 4.567777992104668, 8.899072093526586), (5.064428774391923, 2.3873615305686604, 6.311315303507673), (7.121254328085777, 3.8929371433690307, 6.436047554040005)),
    ((0.012811232785263638, 8.822611491741695, 9.234907083701472), (7.45680438953131, 0.9966169061222518, 7.606829472498982), (9.47976074712619, 6.04668500154162, 6.341579985912633), (3.1368445127260225, 9.719149960716248, 0.2938677471607043), (3.0993985616510464, 8.796570552221512, 4.869520180242636), (3.4931667742298913, 6.618747901270023, 4.016517091011451), (8.027582433935004, 3.695254210546387, 9.599925472912652), (5.058631163489039, 3.244011424562289, 7.463785567090548), (6.9442846245304075, 2.225915273482287, 3.649487804723641), (0.29722902852075683, 2.154388253164475, 7.7915836995422305), (1.4347173832859228, 8.119643333025103, 3.1577523330209276), (2.792764806805735, 0.5491082041895778, 3.210306327006094), (1.778184771364556, 1.024999105969171, 5.171437944957926), (5.101712912933802, 3.7180261324920716, 8.208133764194447), (9.481574778343205, 1.5143794152290813, 6.019147596936579), (8.474533997637733, 1.5991703431401727, 7.491631195223409), (0.4837332607479705, 0.9782095122789713, 7.018530571576946), (0.5158600256550017, 1.7792423554955772, 8.011308041123094), (6.707828665571165, 1.3837125565755426, 4.2807756150793335), (1.0692224170923792, 8.18725827388685, 9.678844004764287), (9.523307677224153, 7.436484057672194, 8.208805537423986), (7.121018451107885, 2.3747961878864032, 6.183922866531483), (3.0353049889069106, 5.130227978364491, 8.265416412204678), (9.383853102547402, 7.988997868097487, 4.316626536280386), (9.861573059745737, 1.367191001555682, 7.771999543109257), (8.89031097513307, 2.261560248844093, 0.1438757134875812), (8.438682977452492, 7.503583421941373, 2.7070165833095605), (0.4149188650710889, 7.195760597330435, 4.795669951751806), (4.550270578371846, 6.465952231246886, 8.40689507897969), (5.3588692823278485, 2.3871962541112257, 4.552941294742845), (5.345384811255986, 1.142337461610211, 0.15719027924801066), (4.670860495161746, 0.8285747932646337, 1.0240855669106474)),
    ((6.145423318805177, 8.469691408207002, 7.264476751683144), (4.794807661770436, 2.8893978293740274, 5.284334371886407), (7.116546434389068, 7.5136529391423625, 4.549582890644704), (5.507671951182871, 3.606937053643462, 0.44130211316144363), (3.057873074732412, 9.48635557827253, 8.683741274514206), (7.284114753707777, 4.636967357208769, 7.191382741817861), (0.801202691328895, 3.2374851286028115, 4.7605677229689745), (5.152525576267806, 8.4148067366799, 3.141191636285383), (4.769985120666782, 2.429610972447377, 5.36188427976358), (4.800116331062451, 5.57345660412857, 7.088318644421925), (9.255441355164203, 4.047473536513026, 8.26086515587658), (8.607522613074853, 0.1489503029663164, 0.5376716454593644), (4.096284474443587, 1.4332165297505017, 2.4072935893230207), (4.868086754118703, 9.943273934485735, 1.3719954568189674), (0.14237450867308543, 3.060720084295838, 2.163802648364672), (3.0869456751459556, 6.365800166782456, 6.251796829113462), (7.931542081409946, 9.411777159322941, 0.34752971174936254), (9.201794556076969, 5.688109668461693, 0.8195675927595303), (6.893772487557755, 8.683746867708033, 3.497459416403663), (8.235276191858492, 6.763703106259561, 2.993395826267027), (2.2579978483045893, 2.9718361977431798, 6.158387685233632), (2.7206100652088114, 0.6664649139484691, 2.1850443978329945), (2.852009987205334, 5.941488697061477, 8.720386083329299), (7.698086292884936, 6.262997760844444, 0.645948622298429), (6.852637208062625, 8.015791187836843, 6.77425768643257), (8.148576815465564, 4.201741573576205, 3.304333925565829), (2.165462204662293, 5.01816524197438, 7.825457277410824), (6.6068261931448005, 7.501072272519407, 7.413007249976262), (1.0643398048148023, 0.44350792804536576, 7.8895153249384755), (0.9581223247580306, 4.69741180022364, 3.8165835763439904), (7.806883191428591, 5.8210274186976605, 5.643692610062194), (5.305695775632394, 5.197332749281436, 3.4573147718660726)),
    ((8.916173265048887, 0.7964832002728928, 9.675734593026245), (6.4506436127281574, 2.398056129224427, 1.9047924901754265), (9.090723221704733, 9.93812066855352, 8.147774494457853), (9.741187475250687, 7.243002898467986, 4.797101633174854), (7.850099530127352, 1.5253108693234674, 4.645938050971693), (6.465997575575874, 8.410339149493101, 5.068767749282444), (9.14491517283752, 6.150863223537877, 9.885859452197229), (2.295922173278705, 7.310715563380431, 9.002977314076874), (4.0463615630295955, 3.1291625059727837, 8.55430667924469), (4.9047047479234065, 6.963134161310542, 3.6025111365401976), (5.672843611720464, 3.203671432457339, 3.8517792574753082), (1.667347872681152, 5.013495945725502, 7.876443779008811), (4.991604288626251, 5.763302730533971, 0.28961108522257417), (2.7873253247604914, 5.733761946138843, 6.81920402206175), (7.821399575246102, 8.340388642092284, 4.901976224994909), (6.51157927514717, 0.800071426544362, 9.091019402963264), (0.7840892436628577, 3.90766745052331, 3.5245129798814254), (2.249603452569515, 7.128413744544114, 7.709819016966191), (5.210720474169854, 3.4394196152666376, 5.303091906400578), (2.2575171492518695, 0.8748124146124514, 7.0328913877824695), (7.474381262306549, 7.514845043501213, 2.399682918292414), (2.212225405599826, 6.7333397313171, 0.39444449174253826), (3.737963122259539, 7.757612977664101, 5.3176829819427915), (4.3522422752508785, 0.7766257028098944, 2.8946429842340047), (0.5525001940055796, 7.280005165185779, 2.9430775336338764), (4.063796811419019, 2.8900739897102854, 1.9943030783608384), (5.93400014689673, 1.2627345972368098, 9.62979378775235), (6.090502012658953, 7.748124719889602, 2.9839020635377587), (0.38914544378182203, 3.7332470998920932, 7.545655369902256), (8.684790483002088, 9.324302727009751, 5.1598958898769585), (8.66961801771549, 3.949483803464796, 1.0966971222943867), (3.119141297448844, 0.2828094310778595, 7.982305449840037)),
    ((5.699140590839665, 6.145218822175122, 2.09251184159939), (2.012294472299666, 8.081716599828814, 4.596840616106062), (8.18934243752212, 6.8826896985583, 9.278941030244548), (9.27982402468389, 4.746930819654075, 0.20049486294124508), (4.2500221182577205, 4.747784593875029, 1.9278908219197022), (0.5717290624334392, 5.0540845739884235, 8.903385334462264), (9.808538273357815, 5.811251274097878, 2.7421221899582005), (6.141680472455274, 5.632203726603221, 5.5780095107460195), (8.262372522882588, 5.2482547348605575, 8.966983607462648), (0.47215665348659397, 3.835251871315213, 8.769911807072992), (5.026105281398946, 1.5136987971663807, 5.880939317117758), (1.1285752485198608, 9.503286157287352, 5.841636223239998), (2.96374690346859, 7.2838183583071086, 7.361034418156941), (4.575092642910269, 0.2578180408731823, 5.118996047385234), (8.934260012934113, 9.81571330625554, 5.7690917566555076), (0.04243922226629171, 9.997580680125564, 8.483218202415726), (2.8022256636343212, 1.4673338862031449, 9.398208149154033), (2.801104053779463, 9.913068982720924, 5.13662431480946), (6.827869725644989, 6.88209949817852, 5.903155373892183), (8.030731324879602, 1.1253233919502936, 1.462431722444698), (5.792140609471063, 2.0124097825901375, 3.2366496698094904), (7.446931136506824, 7.2427023653974345, 0.9984379405938737), (4.962420445130881, 6.880940233734188, 9.919554727528467), (1.6853629385739888, 9.145027056032747, 2.711910143817544), (3.5241276335540404, 1.8578147172298676, 2.62392092010445), (7.748781433301759, 2.50498078589634, 4.148353563197462), (9.229644036370704, 6.551213360027881, 4.578360683025407), (3.4366170898505635, 1.6446578912739818, 1.8989276067836869), (4.147385525730486, 2.067966421964784, 3.0397338416904205), (9.461622460292386, 2.359655076606597, 0.1944900782137038), (2.446574878656036, 9.572016544918498, 8.511011413581889), (0.0049885181571718284, 7.4713199316620145, 4.494037590176042)),
    ((6.244046142458906, 2.9614632789929485, 1.042473346106303), (6.124532045401484, 0.8197190164872337, 6.342770842936392), (0.673582770670248, 2.3565161345911934, 9.892665599462688), (9.804958639537983, 6.999361666144015, 8.421299328736854), (5.109856727564466, 9.454913067425135, 7.139040975690395), (1.9231109070725283, 4.673195398037206, 5.99515898381213), (9.813172900629555, 2.929795260397039, 7.301312992023558), (6.858715575101009, 8.76097699795155, 4.153828953415195), (8.151603981860983, 9.927360151733593, 3.0223190140931133), (0.03650371105003658, 3.9474506099516526, 6.735972419309734), (5.27107876925224, 3.7759956055159414, 5.169919166365854), (3.5389492093484733, 6.647156743178804, 3.8375840122659466), (8.91003675950515, 7.747714119494187, 5.737029922766426), (9.76977584825002, 2.161619776674748, 7.429697088514352), (8.126522920473093, 7.114724108850938, 5.216582185300725), (2.539773370005889, 1.5539191279743825, 4.571167402525593), (4.454140932988566, 6.606717021588811, 5.903189128597337), (3.3767778681338303, 6.165254873191603, 1.4381915254729893), (9.31559651712774, 9.639554393365966, 7.0626848654066645), (0.4870867450788363, 8.052121057926096, 9.858707429733464), (1.75587684183653, 3.480215144062495, 1.6598510409834621), (1.4543382736494082, 3.7443722497737153, 4.927340652408124), (3.520659891435457, 8.636530337870422, 4.174661640771397), (4.85868271016924, 5.365046011714077, 4.5808038694344155), (2.0049356227417094, 2.1043087727864673, 4.215592157159968), (3.791216955717357, 4.1174052145822415, 4.90708426091528), (7.668676519263845, 5.542871835828498, 2.514258269209808), (5.840883354893414, 8.862656372466745, 1.2284806914422264), (0.5870778100736085, 6.0704127386593925, 9.498144984191317), (1.4539230211233767, 0.12709657926542106, 8.04848627666273), (2.748242533313902, 9.293751305221209, 0.3830581513835307), (4.156871656592607, 4.8428306146019775, 6.239622769867239)),
    ((1.3222875477886387, 5.819447677115754, 3.8769458906164402), (8.788973844201802, 3.007203443941088, 8.149668781613807), (7.315225495197919, 0.3824076625261408, 2.314958748602154), (5.931810329937651, 9.649865851645007, 2.1880971659802873), (6.084477483927233, 5.574748390850301, 3.3467738462205032), (1.1943992473493203, 2.8559472629867, 4.856095761320088), (7.168491874590836, 0.7743259454734241, 2.0800339296883252), (0.19520000216485922, 9.601812208452923, 5.0169303013551305), (9.787216109037118, 3.471590060708337, 1.2661039217210912), (0.5630096497153358, 7.52338513012226, 7.112886200873469), (0.8211787372139179, 4.578384994411734, 0.8433739171875176), (7.235544400219042, 3.5630290161469027, 8.736986401480477), (7.0146658783071185, 7.239630152072976, 2.5602483636071813), (3.8707277756680245, 8.421683603831173, 0.400391131020128), (5.635251918226237, 8.443126190711407, 4.563163153675718), (9.882559366465438, 0.6298021896190475, 8.950938639921844), (8.839205778016906, 1.3998992939674249, 6.207121539707239), (4.526492947250206, 4.469938213672128, 4.863187865836146), (1.5817723519234395, 7.134468190317767, 1.8419406918441417), (5.66154049817284, 7.134904237778658, 1.6020996190273051), (9.6638054861471, 4.740523589283798, 9.791682508212197), (9.30125081823199, 7.132125288716812, 7.4064570224560065), (9.788731474116814, 2.1535825548983856, 2.664796265775257), (9.26510977986367, 1.6058667516375014, 8.246878706861587), (8.272619878066525, 1.8173837618967215, 5.282638291226119), (2.3054117980589406, 1.0389666756217952, 3.12930111233337), (4.047534697405486, 6.364842999993009, 0.5120254412006953), (4.916305260014065, 3.094185114440929, 9.571410342352497), (8.682314031197595, 4.760354425878561, 7.106211136408815), (0.1720900589513752, 4.295846567470862, 7.4099157341684), (0.4034430417439816, 8.081948780362502, 7.551538755468666), (3.080594255131466, 0.8274623924482805, 3.8069731233191617)),
    ((4.382260819508446, 3.5845360584396477, 4.509500019832247), (2.588033543208035, 4.651435602980389, 9.832612322792016), (6.00036283187023, 2.646767384117117, 3.589875512987918), (5.852359882925892, 6.0196333692904656, 1.4930859582413214), (3.701654012840395, 7.613917214717333, 3.300784842123534), (0.05320814587702727, 4.138779674655597, 3.7825495859577973), (7.585687762329398, 2.0209781700204665, 5.106394922033642), (6.55138282106773, 2.21423046005771, 1.5820325968112048), (3.473063304248888, 5.251393643215721, 9.330544618993802), (9.073915554180306, 0.7211337342735891, 2.277556960916718), (7.518250092878222, 0.30832490717524696, 9.460532200135189), (0.22475080056905128, 0.6108516361866589, 5.113716020044896), (0.47676021054967155, 7.2495051826864385, 6.530774688213255), (7.250815230902921, 9.48254140036942, 5.9921271699013525), (7.92216719461721, 3.227975524061896, 3.0399709652677522), (3.102925824985854, 2.9865980315153573, 6.437340908759424), (2.3648297075315927, 3.1617967773599442, 5.531733288555481), (7.6172079210847965, 8.258189133116883, 8.706433481133574), (3.0385395418950747, 9.231866786531086, 6.441522112769315), (1.4736575137554753, 5.379503628337318, 7.835359514889025), (9.794309170659997, 5.327269941611691, 5.162949149398748), (0.40156135617521627, 4.108398399306576, 2.571461005037806), (3.9757614913135484, 6.8848144134749685, 3.858916735090774), (1.5069706908205538, 9.876316271945045, 5.467731109709238), (3.6032410613649968, 1.8941633195362895, 5.133340115101458), (3.150909462536559, 8.219700755858378, 4.366981754148522), (3.6569722395743964, 0.6558584830422831, 0.8405720105278125), (6.31863636970436, 3.2623478440360287, 4.922260359215864), (5.430007959437736, 9.393618348416696, 1.245520310340098), (0.1613567423476081, 9.75620311545086, 6.201998377575469), (1.2224970646318623, 4.9245314663497055, 3.82965358193513), (4.115186274072091, 8.500938778826136, 8.083709865196958))
    );    
 
constant k_height  : integer := 3;
constant k_width   : integer := 3;
constant k_depth   : integer := 3;
constant k_filters : integer := 16; 

constant kernel : float_4d_vector :=
    (
    (((7.025540099322349, 8.286202573468106, 9.886344144646898, 0.10268289160940247, 9.369615907788685, 4.1247207350372825, 8.3037461331318, 8.89039029586693, 4.618194622665448, 8.185996583234132, 7.742818419413451, 9.577505066390735, 3.9864302165035035, 8.907562360305242, 6.289454305067439, 8.56476307603003), (4.577210520507507, 0.20040252717530405, 5.103757955207136, 8.059229643889875, 8.070645390035374, 4.477810848128879, 1.1483696517707964, 0.8729833057055125, 6.749685221232817, 9.477900976739665, 9.840827793951835, 6.598919388020108, 9.577377603091769, 1.4235206725739458, 8.727515788376085, 9.926462202168665), (0.18035469413071326, 0.7507892446350917, 0.15239097114680633, 3.6582770774991302, 4.32471338469325, 2.4836168204097864, 8.925153530820536, 5.858635678931959, 9.393379149453322, 5.660233562615197, 6.143951046877552, 1.824748722376699, 6.16990798242532, 8.025216218842422, 3.075365261468148, 5.691569462461485)),
    ((0.5908512535629828, 1.9414928755523786, 5.304067938060132, 0.012636501553888735, 0.20704119218057593, 0.3375596272844339, 6.819274293782422, 4.266702351764443, 5.0036941130220995, 8.580123382403539, 2.0245483959921264, 3.4294057411653833, 4.391852981463264, 6.0548679657589135, 2.968222529361592, 3.7505796956213935), (8.328898882479592, 8.053656054031128, 9.758883762934706, 0.28216093019822197, 0.9032945489967414, 3.035847352895394, 1.99597969311486, 5.664972373455016, 1.4388362913684283, 0.8550254589272022, 7.729183197876075, 0.13983082356815446, 8.456352779869219, 8.66643219957237, 8.953603236493574, 9.681609869192368), (1.766465333165762, 5.153729397640269, 9.670715341761797, 0.38455878259616827, 5.0110722591849735, 8.192810946324805, 0.294276364736179, 3.6917642067585312, 0.6181400388582936, 5.405621769701133, 9.617404382706324, 3.4283799846497107, 5.765581646682662, 6.606387937914711, 4.777651397950194, 3.3111467645002826)),
    ((5.522414563993685, 7.866642961885636, 4.783342787514417, 2.9971781484111846, 6.896770735283148, 4.5363575923391934, 8.006685226208102, 1.1264889601501427, 2.0630195731894494, 9.360688511594196, 2.646372419329021, 9.744908756531936, 4.815026076271231, 5.965257469789968, 8.741682885257948, 8.209903797313054), (1.6768976129965174, 1.2189973564761725, 3.8773191373923277, 5.097582158423339, 1.9093706655215237, 8.488432820981378, 3.8003635507069413, 2.168311810358121, 0.7489458105308078, 1.06089971874895, 4.0929736971679445, 3.039810920394749, 0.8933915793718916, 1.0203220218201625, 7.188369634522265, 8.66428596343897), (1.2652483098095912, 7.886088536706319, 7.766146752671281, 8.284710157544264, 0.7496031454734964, 6.076967904539065, 7.610417309848904, 5.689609451340734, 0.8787596567551226, 2.0738110138011603, 7.580691843252368, 1.9054830448495474, 3.2770838270698244, 6.042348214576889, 9.791162399465552, 5.47899743260316))),
        (((5.34886000092981, 1.7287064375285555, 8.294613412436759, 4.394378149140191, 7.42960074478529, 2.7974304084351242, 4.965402336579175, 7.36304316765807, 4.74993557609002, 1.3721884553465824, 9.694519585971385, 6.615226014346628, 8.950403563602826, 8.459517168568807, 8.85036515193919, 0.8307004482573244), (7.334328555939074, 8.974945002048624, 6.655507260366232, 1.6998276526267697, 8.412191501407635, 8.303721565482308, 7.10302256566205, 3.823697062772525, 4.550239958920102, 8.978409947819078, 0.9905189061648079, 1.3871178919831273, 8.75264221586211, 7.460225608269814, 3.133395267744344, 7.055351772923576), (7.986683770597475, 9.863580888159726, 4.267429829715858, 5.357092620665082, 8.991369306753322, 5.015281532425034, 1.316239212468736, 4.423734972525542, 8.022603918014127, 8.305410291712567, 0.05395725599876222, 2.9959520578074503, 8.246124226316503, 4.964701253213923, 1.2793917000963628, 4.124660944174888)),
    ((4.348145201683514, 8.491919970618953, 3.179640110669686, 5.60227103873463, 9.643180988071158, 1.4133748250074707, 4.177102263564741, 7.654738692556517, 0.8392787787981049, 6.843714897905517, 0.3426965172406804, 8.572838441680808, 9.403944856969913, 7.510544016773155, 9.408651585416141, 6.645714779762511), (9.393837735974467, 9.329119747066105, 7.307381944800375, 1.556089219835467, 8.669958175114015, 4.532442908291269, 6.55341464922821, 8.86719076140458, 0.09612078256113987, 3.3464403368480733, 0.11586458584766146, 5.790010597886923, 2.768352894535926, 0.5316243714671309, 6.445056099286344, 2.054130893707913), (2.057679948774979, 8.28713063531413, 0.9920479825526429, 7.652729959640785, 6.820987882812371, 1.7246232616170865, 3.893666547885851, 4.019780798420021, 3.0501165611497005, 6.550005514457297, 4.7563889594226545, 4.317803312116803, 3.414217769941481, 7.73039305447479, 5.145235183612971, 8.010909148210082)),
    ((7.1369560652159505, 9.819140462635257, 9.709277745228546, 7.997091783482255, 0.7334475914347449, 5.851919122006431, 5.079728325429357, 5.592874934708157, 3.1091064790731693, 9.255957500076239, 8.806358926817682, 3.7390581023821667, 5.281486161893508, 1.9585282362938106, 8.410495017303893, 4.814839059887105), (1.8924215589580018, 9.49191358354193, 2.86017570678631, 1.2450122594871793, 5.484864661156358, 5.322775684253717, 8.587525990395623, 3.0590255391122545, 4.471762845577727, 5.479935334939451, 7.955406641228571, 6.5922359880375625, 1.0932190136053854, 2.098164619219114, 1.5959318958319868, 2.4087597421609495), (3.9346415917414044, 4.36836932275817, 5.671464232070757, 6.820937905783801, 1.0200556798974492, 9.909677059237493, 9.835972975087673, 1.8728678222283557, 9.79021435966103, 1.3036519212043862, 4.386122931343842, 6.02788950835245, 2.988613318776119, 8.727409747718104, 0.166210370581803, 1.9297599977343982))),
        (((1.0758925002103858, 7.70676422347084, 8.692085218032647, 2.648825469173092, 1.5072698748157942, 7.094061677730749, 8.456226718694762, 5.517466256097336, 4.637590126389268, 7.144232030083668, 6.6787176332717335, 2.3684722167083585, 6.085533576370807, 8.693062429188258, 4.549495249287223, 6.189829573933633), (1.2172759554816837, 9.703711206508938, 7.894585128058741, 8.916707751754585, 2.2734540548299975, 7.861100857834721, 3.902910165989426, 4.163898192200967, 0.17402818520258712, 3.700067095175884, 0.014014409380317394, 2.0200810929316404, 8.960315859473617, 1.1919964348551593, 0.8961621031795908, 1.521951944155281), (7.225274638507308, 9.097435234855032, 8.873137599530423, 9.184413131994875, 2.189177235808706, 7.313898067673633, 0.7279770188497803, 6.640937671075406, 6.019325455343418, 6.997360354153001, 5.1914956445052525, 3.4540115826429174, 6.677806159136517, 5.375769788921735, 6.378118150449742, 2.8989214698302304)),
    ((9.947798987258562, 0.13382257467489334, 6.711680152596255, 6.152768360313657, 3.882275520386118, 3.6689079227214503, 9.139092093640972, 8.114894721921983, 5.818499758991509, 4.5494433117244935, 8.18029387251931, 6.019490065007739, 0.49997523826237233, 6.238117115150182, 5.373579057671344, 3.6175359900146464), (6.029996687899729, 3.980359154279003, 6.650848881050324, 3.1305066331195386, 0.40335499154453003, 2.989432652961569, 0.07084825520495608, 8.367492478388918, 5.414041476100996, 4.676696605008123, 1.321301570663681, 5.685525156914332, 4.575451254199983, 9.661020841678873, 0.7558110411170749, 2.867697021031627), (3.3888725000986497, 2.45058717623331, 4.5623421982215, 1.2173360149441637, 7.393978810449898, 4.492541064995833, 1.6346216220170318, 2.9965397670310834, 3.8255119219797074, 7.9298707426315, 5.019017724738375, 1.1485317884526514, 4.4442778285264914, 4.459910761478595, 4.497284605286559, 5.368692623505266)),
    ((4.7112217353960775, 9.399275210242747, 8.987435862036408, 8.183107965243137, 7.30368992975065, 1.1592570750178488, 1.2686097607865976, 5.457730548859304, 9.511432150611533, 6.527126018079796, 1.9438544749145792, 4.153273334325687, 2.516991137087908, 9.41362906520949, 6.1797311907555, 9.837347794937656), (9.651717514837033, 0.9843587131255938, 6.85714488174094, 1.23377586223555, 0.8387158712310228, 1.9015907440344737, 6.875051725078475, 0.03415151503306846, 3.6046349976209657, 5.5107894001610696, 5.453775019661965, 1.7329898783877895, 3.439466591559348, 9.3770726446942, 4.059278464384378, 7.968339668387763), (4.599364435742629, 1.5543104490667692, 3.0439107010643807, 2.2319049574826924, 6.073580111401759, 3.529961821663382, 9.598158524504845, 4.492132490942552, 1.9486329544675063, 8.249232889467633, 8.523554941562756, 9.053601629043934, 0.977642836407564, 0.9694329982534899, 1.3146138388569828, 3.6209752579179355)))
    );
 
constant gamma : float_1d_vector := 
    (
    3.2638158798217773,
    4.460397720336914,
    1.18198561668396,
    1.6533160209655762,
    4.321843147277832,
    1.6785709857940674,
    4.001209259033203,
    6.566650390625,
    2.339569568634033,
    3.654820442199707,
    3.554124116897583,
    3.6159822940826416,
    2.8188273906707764,
    2.1044859886169434,
    3.7799949645996094,
    1.9643325805664062
    );
constant beta : float_1d_vector := 
    (
    -2.890369415283203,
    -6.697666645050049,
    0.5552693009376526,
    0.7817191481590271,
    -4.420159339904785,
    0.9831221699714661,
    -4.607707500457764,
    -9.767300605773926,
    -0.3404657244682312,
    1.0352110862731934,
    0.7899404764175415,
    0.9098617434501648,
    0.32240909337997437,
    -0.10215473920106888,
    1.3165702819824219,
    1.1973998546600342
    ); 
constant moving_mean : float_1d_vector := 
    (
    -0.7467830181121826,
    0.406264990568161,
    0.058190274983644485,
    0.06197834387421608,
    -0.036936476826667786,
    -0.0039504277519881725,
    -0.03281150385737419,
    -1.057032823562622,
    -0.03209839388728142,
    0.043669186532497406,
    -0.0017793704755604267,
    0.05360546335577965,
    -0.23466050624847412,
    -0.00626344932243228,
    0.017854779958724976,
    -0.1660752296447754
    );    
constant moving_variance : float_1d_vector := 
    (
    0.1594277024269104,
    0.04255719110369682,
    0.19109822809696198,
    0.4208472967147827,
    0.14984990656375885,
    0.013252475298941135,
    0.12210448086261749,
    0.2738870084285736,
    0.059880033135414124,
    0.7717112898826599,
    0.6764482855796814,
    0.8243041038513184,
    0.3935566246509552,
    0.1252153068780899,
    0.7929491400718689,
    0.37377357482910156
    );        
   
 constant epsilon : real := 0.001;   
    
BEGIN       
    process (CLK, reset)
        
    -- kernels variables
    variable n_i_height : integer := (i_height - k_height) + 1; 
    variable n_i_width  : integer  := (i_width - k_width) + 1; 
    variable n_i_depth  : integer  := (i_depth - k_depth) + 1; 
    variable conv_sum   : real := 0.0;
    
    -- imgage variables
    variable temp_img  : float_3d_vector (0 to (n_i_height - 1), 0 to (n_i_width - 1), 0 to (i_filters - 1)) := (others => (others => (others => 0.0)));
    
    -- batch norm variables
    variable x : real := 0.0;
    variable x_norm : real := 0.0;
    variable y : real := 0.0;
    
    -- activation variables
    variable act_x : real := 0.0;
    
    -- max pool variables
    variable max_val : real := 0.0;
    variable mh : integer := 0;
    variable mw : integer := 0;
    
    begin
        if reset ='1' then                          
        elsif(CLK'event and CLK='1') then
                                  
            -- perform conv
            for d in 0 to (n_i_depth - 1) loop -- performed only once
                for h in 0 to (n_i_height - 1) loop
                    for w in 0 to (n_i_width - 1) loop
                        for k_f in 0 to (k_filters - 1) loop
                            conv_sum := 0.0;
                            for k_d in 0 to (k_depth - 1) loop
                                for k_h in 0 to (k_height - 1) loop
                                    for k_w in 0 to (k_width - 1) loop
                                        conv_sum := conv_sum + img((h+ k_h), (w + k_w), (d + k_d)) * kernel(k_h, k_w, k_d, k_f);
                                    end loop;
                                end loop;
                             temp_img(h,w,k_f) := conv_sum;   
                             end loop;            
                        end loop;
                    end loop;
                 end loop;
            end loop;            
            
            -- perform batchNorm 
            for h in 0 to (n_i_height - 1) loop
                for w in 0 to (n_i_width -1) loop
                    for d in 0 to (k_filters - 1) loop
                        x := temp_img(h,w,d);
                        x_norm := (x - moving_mean(d)) / ((moving_variance(d) - epsilon) ** 0.5);
                        y := (gamma(d) * x_norm) + beta(d);
                        temp_img(h, w, d) := y;
                    end loop;  
                end loop;
            end loop;
            
            -- perform LeakyReLU
            for h in 0 to (n_i_height - 1) loop
                for w in 0 to (n_i_width -1) loop
                    for d in 0 to (k_filters - 1) loop
                        act_x := temp_img(h, w, d);
                        if (act_x > 0.0) then
                            temp_img(h, w, d) := act_x;
                        else
                            temp_img(h, w, d) := -0.01 * act_x;    
                        end if;     
                    end loop;  
                end loop;
            end loop;
            
            -- perform MaxPool
            for d in 0 to (k_filters - 1) loop
                mh := 0;
                for mh_outer in 0 to ((n_i_height - 2) / stride) loop
                    mw := 0;
                    for mw_outer in 0 to ((n_i_width - 2) / stride) loop
                        max_val := temp_img(mh, mw, d);
                        if (temp_img(mh, mw + 1, d) > max_val) then
                            max_val := temp_img(mh, mw + 1, d);
                        end if;
                        if (temp_img(mh + 1, mw, d) > max_val) then
                            max_val := temp_img(mh + 1, mw, d);
                        end if;
                        if (temp_img(mh + 1, mw + 1, d) > max_val) then
                            max_val := temp_img(mh + 1, mw + 1, d);
                        end if;
            
                        new_img(mh_outer, mw_outer, d) <= max_val;
            
                        mw := mw + stride;
                    end loop;
                    mh := mh + stride;
                end loop;
            end loop;

        end if;
    end process;
end Behavioral; 
